// I should wite example top_here here 