// I should wite example tb here 