// I should wite example base_test here 